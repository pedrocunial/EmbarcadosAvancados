
module niosHello (
	butaos_export,
	clk_clk,
	reset_reset_n,
	leds_1_name);	

	input	[4:0]	butaos_export;
	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	leds_1_name;
endmodule
