
module niosHello (
	butaos_export,
	clk_clk,
	leds_1_name,
	reset_reset_n);	

	input	[4:0]	butaos_export;
	input		clk_clk;
	output	[3:0]	leds_1_name;
	input		reset_reset_n;
endmodule
